import p_alu::*;

module m_alu(
	input s_control control,
	output[31:0] result,
	output e_cmp_res cmp_res
);
endmodule