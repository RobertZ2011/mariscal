module m_control;
    
endmodule