`timescale 1 ns/10 ps

module decoder_test;
    initial begin
        $finish;
    end
endmodule